module led_driver(

);
endmodule
